// Types.bsv
// 공통 타입 정의 및 인터페이스

package Types;

// 기본 타입 정의
typedef 64  TIMESTAMP_WIDTH; // Unix timestamp 비트 폭

endpackage